/* 
    Author          : Abhinav Nandwani
    Filename        : CommTB.sv
    Description     : This module is a testbench for the 
                      RemoteComm.sv and UART_wrapper.sv modules.
*/

module CommTB();

    
