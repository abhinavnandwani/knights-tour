module SPI_mnrch_tb();


    























endmodule